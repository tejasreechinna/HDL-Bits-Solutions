module top_module( input in, output out );
wire x ;
    assign x=in ;
    assign out=x;
endmodule
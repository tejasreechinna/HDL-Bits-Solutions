module top_module (
    input in,
    output out);
 wire w ;
    assign w=in;
    assign out=w;
endmodule

module top_module ( input a, input b, output out );
    mod_a dut (a , b , out);
endmodule
